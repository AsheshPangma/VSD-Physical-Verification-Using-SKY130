magic
tech sky130A
timestamp 1665494037
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628528476
transform 1 0 230 0 1 0
box -19 -24 65 296
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665494037
transform 1 0 0 0 1 0
box -19 -24 249 296
<< end >>
