* NGSPICE file created from inverter.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_RV7F6E a_n173_n150# a_n78_n150# a_63_n238# a_n129_n238#
+ w_n311_n360# a_114_n150# a_18_n150# a_n33_172#
X0 a_114_n150# a_63_n238# a_18_n150# w_n311_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=180000u
X1 a_n78_n150# a_n129_n238# a_n173_n150# w_n311_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=180000u
X2 a_18_n150# a_n33_172# a_n78_n150# w_n311_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=180000u
C0 a_114_n150# a_n173_n150# 0.05fF
C1 a_n33_172# a_63_n238# 0.02fF
C2 a_n33_172# a_n78_n150# 0.00fF
C3 a_114_n150# a_18_n150# 0.23fF
C4 a_n173_n150# a_n78_n150# 0.23fF
C5 a_63_n238# a_18_n150# 0.00fF
C6 a_n33_172# a_18_n150# 0.01fF
C7 a_18_n150# a_n78_n150# 0.23fF
C8 a_63_n238# a_n129_n238# 0.04fF
C9 a_n33_172# a_n129_n238# 0.02fF
C10 a_n129_n238# a_n78_n150# 0.00fF
C11 a_18_n150# a_n173_n150# 0.11fF
C12 a_n129_n238# a_n173_n150# 0.00fF
C13 a_63_n238# a_114_n150# 0.00fF
C14 a_114_n150# a_n78_n150# 0.11fF
C15 a_114_n150# w_n311_n360# 0.19fF
C16 a_18_n150# w_n311_n360# 0.13fF
C17 a_n78_n150# w_n311_n360# 0.13fF
C18 a_n173_n150# w_n311_n360# 0.19fF
C19 a_63_n238# w_n311_n360# 0.21fF
C20 a_n129_n238# w_n311_n360# 0.21fF
C21 a_n33_172# w_n311_n360# 0.16fF
.ends

.subckt sky130_fd_pr__pfet_01v8_6LLYWG VSUBS a_n33_131# w_n311_n319# a_114_n100# a_63_n197#
+ a_18_n100# a_n129_n197# a_n173_n100# a_n78_n100#
X0 a_18_n100# a_n33_131# a_n78_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 a_114_n100# a_63_n197# a_18_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X2 a_n78_n100# a_n129_n197# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
C0 a_n78_n100# a_114_n100# 0.07fF
C1 a_18_n100# a_n78_n100# 0.16fF
C2 a_n78_n100# a_n129_n197# 0.00fF
C3 a_n33_131# a_63_n197# 0.02fF
C4 a_n78_n100# a_n173_n100# 0.16fF
C5 a_n78_n100# w_n311_n319# 0.09fF
C6 a_114_n100# a_63_n197# 0.00fF
C7 a_18_n100# a_n33_131# 0.00fF
C8 a_n33_131# a_n129_n197# 0.02fF
C9 a_18_n100# a_63_n197# 0.00fF
C10 a_n129_n197# a_63_n197# 0.04fF
C11 a_n33_131# w_n311_n319# 0.09fF
C12 w_n311_n319# a_63_n197# 0.06fF
C13 a_18_n100# a_114_n100# 0.16fF
C14 a_n173_n100# a_114_n100# 0.04fF
C15 a_18_n100# a_n173_n100# 0.07fF
C16 a_n173_n100# a_n129_n197# 0.00fF
C17 w_n311_n319# a_114_n100# 0.13fF
C18 a_18_n100# w_n311_n319# 0.09fF
C19 w_n311_n319# a_n129_n197# 0.06fF
C20 w_n311_n319# a_n173_n100# 0.13fF
C21 a_n33_131# a_n78_n100# 0.00fF
C22 a_114_n100# VSUBS 0.01fF
C23 a_18_n100# VSUBS 0.01fF
C24 a_n78_n100# VSUBS 0.01fF
C25 a_n173_n100# VSUBS 0.01fF
C26 a_63_n197# VSUBS 0.13fF
C27 a_n129_n197# VSUBS 0.13fF
C28 a_n33_131# VSUBS 0.13fF
C29 w_n311_n319# VSUBS 2.53fF
.ends

.subckt inverter in out vss vdd
XXM1 out XM1/a_n78_n150# in in vss XM1/a_114_n150# out in sky130_fd_pr__nfet_01v8_RV7F6E
XXM2 vss in vdd XM2/a_114_n100# in vdd in vdd XM2/a_n78_n100# sky130_fd_pr__pfet_01v8_6LLYWG
C0 vdd in 0.97fF
C1 out in 0.77fF
C2 XM1/a_n78_n150# out 0.12fF
C3 XM1/a_114_n150# in 0.00fF
C4 vdd XM2/a_n78_n100# 0.12fF
C5 out XM2/a_n78_n100# 0.12fF
C6 XM1/a_n78_n150# in 0.06fF
C7 vdd out 0.29fF
C8 XM1/a_114_n150# out 0.12fF
C9 XM2/a_114_n100# vdd 0.12fF
C10 XM2/a_114_n100# out 0.12fF
C11 XM2/a_n78_n100# in 0.06fF
C12 XM2/a_114_n100# vss 0.01fF
C13 XM2/a_n78_n100# vss 0.01fF
C14 vdd vss 3.51fF
C15 in vss 2.52fF
C16 XM1/a_114_n150# vss 0.32fF
C17 XM1/a_n78_n150# vss 0.26fF
C18 out vss -1.81fF
.ends

