magic
tech sky130A
magscale 1 2
timestamp 1665423701
<< pwell >>
rect -58 646 569 1267
rect -60 645 569 646
<< metal1 >>
rect 148 2390 348 2528
rect -48 2018 592 2390
rect -112 1936 290 1982
rect -112 1652 -56 1936
rect 534 1898 592 2018
rect 94 1868 592 1898
rect 189 1684 616 1718
rect 552 1678 616 1684
rect -112 1604 384 1652
rect -538 1416 -338 1474
rect -112 1416 -56 1604
rect -538 1360 -56 1416
rect -538 1274 -338 1360
rect -112 1142 -56 1360
rect 554 1440 616 1678
rect 816 1440 1016 1498
rect 554 1368 1016 1440
rect -112 1086 294 1142
rect -112 726 -56 1086
rect 554 1048 616 1368
rect 816 1298 1016 1368
rect 94 1008 616 1048
rect 190 782 598 806
rect 190 762 600 782
rect -112 670 384 726
rect 486 642 600 762
rect -58 310 600 642
rect -58 308 566 310
rect 144 186 344 308
use sky130_fd_pr__nfet_01v8_RV7F6E  XM1
timestamp 1665423701
transform 1 0 258 0 1 907
box -311 -360 311 360
use sky130_fd_pr__pfet_01v8_6LLYWG  XM2
timestamp 1665423701
transform 1 0 263 0 1 1793
box -311 -319 311 319
<< labels >>
flabel metal1 -538 1274 -338 1474 0 FreeSans 256 0 0 0 in
port 0 nsew
flabel metal1 816 1298 1016 1498 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 144 186 344 386 0 FreeSans 256 0 0 0 vss
port 2 nsew
flabel metal1 148 2328 348 2528 0 FreeSans 256 0 0 0 vdd
port 3 nsew
<< end >>
