magic
tech sky130A
timestamp 1665478438
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1665478438
transform 1 0 0 0 1 0
box -19 -24 249 296
<< end >>
